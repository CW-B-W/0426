wire [15:0] FIR_C [99:0];
assign FIR_C[0] = 16'h1000;    // 1.00000000000000000000
assign FIR_C[1] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[2] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[3] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[4] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[5] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[6] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[7] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[8] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[9] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[10] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[11] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[12] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[13] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[14] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[15] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[16] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[17] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[18] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[19] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[20] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[21] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[22] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[23] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[24] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[25] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[26] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[27] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[28] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[29] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[30] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[31] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[32] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[33] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[34] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[35] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[36] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[37] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[38] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[39] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[40] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[41] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[42] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[43] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[44] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[45] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[46] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[47] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[48] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[49] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[50] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[51] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[52] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[53] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[54] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[55] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[56] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[57] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[58] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[59] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[60] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[61] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[62] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[63] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[64] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[65] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[66] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[67] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[68] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[69] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[70] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[71] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[72] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[73] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[74] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[75] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[76] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[77] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[78] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[79] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[80] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[81] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[82] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[83] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[84] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[85] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[86] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[87] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[88] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[89] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[90] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[91] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[92] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[93] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[94] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[95] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[96] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[97] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[98] = 16'h0000;    // 0.00000000000000000000
assign FIR_C[99] = 16'h1000;    // 1.00000000000000000000
